** sch_path: /foss/designs/real/inyeon-4-chipaton-2025/lvs/gf180mcu_osu_sc_gp9t3v3__maj3.sch
.subckt gf180mcu_osu_sc_gp9t3v3__maj3 VDD VSS A B C Y
*.PININFO VDD:B VSS:B A:I B:I C:I Y:O
XM1 net1 C VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM2 X B net1 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM3 net6 A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM5 net2 A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM6 X C net2 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM4 X B net6 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM7 X B net5 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM8 net5 C VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM9 X B net4 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM10 net4 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM11 X C net3 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM12 net3 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM13 Y X VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM14 Y X VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM15 Y X VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM16 Y X VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
.ends
