magic
tech gf180mcuD
magscale 1 10
timestamp 1753235859
<< nwell >>
rect -145 362 1724 963
<< pwell >>
rect -145 264 1557 362
rect -145 0 1550 264
rect -145 -240 1557 0
<< nmos >>
rect 86 0 206 264
rect 310 0 430 264
rect 534 0 654 264
rect 758 0 878 264
rect 982 0 1102 264
rect 1206 0 1326 264
rect 1430 0 1550 264
<< pmos >>
rect 86 504 186 870
rect 310 504 410 870
rect 534 504 634 870
rect 758 504 858 870
rect 982 504 1082 870
rect 1206 504 1306 870
rect 1430 504 1530 870
<< ndiff >>
rect -2 236 86 264
rect -2 96 11 236
rect 57 96 86 236
rect -2 0 86 96
rect 206 0 310 264
rect 430 142 534 264
rect 430 96 459 142
rect 505 96 534 142
rect 430 0 534 96
rect 654 0 758 264
rect 878 236 982 264
rect 878 96 907 236
rect 953 96 982 236
rect 878 0 982 96
rect 1102 0 1206 264
rect 1326 236 1430 264
rect 1326 96 1355 236
rect 1401 96 1430 236
rect 1326 0 1430 96
rect 1550 237 1638 264
rect 1550 97 1579 237
rect 1625 97 1638 237
rect 1550 0 1638 97
<< pdiff >>
rect -2 816 86 870
rect -3 792 86 816
rect -3 752 11 792
rect -2 652 11 752
rect 57 652 86 792
rect -2 504 86 652
rect 186 504 310 870
rect 410 792 534 870
rect 410 652 459 792
rect 505 652 534 792
rect 410 504 534 652
rect 634 504 758 870
rect 858 792 982 870
rect 858 652 907 792
rect 953 652 982 792
rect 858 504 982 652
rect 1082 504 1206 870
rect 1306 792 1430 870
rect 1306 652 1355 792
rect 1401 652 1430 792
rect 1306 504 1430 652
rect 1530 793 1638 870
rect 1530 653 1579 793
rect 1625 653 1638 793
rect 1530 504 1638 653
<< ndiffc >>
rect 11 96 57 236
rect 459 96 505 142
rect 907 96 953 236
rect 1355 96 1401 236
rect 1579 97 1625 237
<< pdiffc >>
rect 11 652 57 792
rect 459 652 505 792
rect 907 652 953 792
rect 1355 652 1401 792
rect 1579 653 1625 793
<< polysilicon >>
rect 86 962 1306 1022
rect 86 870 186 962
rect 310 870 410 914
rect 534 870 634 914
rect 758 870 858 914
rect 982 870 1082 914
rect 1206 870 1306 962
rect 1430 870 1530 914
rect 86 458 186 504
rect 310 458 410 504
rect 534 458 634 504
rect 758 458 858 504
rect 982 458 1082 504
rect 1206 458 1306 504
rect 1430 458 1530 504
rect 86 264 206 458
rect 310 414 430 458
rect 534 414 654 458
rect 310 401 654 414
rect 310 355 459 401
rect 505 355 654 401
rect 310 342 654 355
rect 310 264 430 342
rect 534 264 654 342
rect 758 414 878 458
rect 982 414 1102 458
rect 758 401 1102 414
rect 758 355 907 401
rect 953 355 1102 401
rect 758 342 1102 355
rect 758 264 878 342
rect 982 264 1102 342
rect 1206 401 1326 458
rect 1206 355 1243 401
rect 1289 355 1326 401
rect 1206 264 1326 355
rect 1430 401 1550 458
rect 1430 355 1467 401
rect 1513 355 1550 401
rect 1430 264 1550 355
rect 86 -92 206 0
rect 310 -44 430 0
rect 534 -44 654 0
rect 758 -44 878 0
rect 982 -44 1102 0
rect 1206 -92 1326 0
rect 86 -152 1326 -92
rect 1430 -152 1550 0
<< polycontact >>
rect 459 355 505 401
rect 907 355 953 401
rect 1243 355 1289 401
rect 1467 355 1513 401
<< metal1 >>
rect -2 849 1414 1029
rect 11 792 57 803
rect 11 264 57 652
rect 459 792 505 849
rect 459 641 505 652
rect 907 792 953 803
rect 1355 792 1401 849
rect 907 606 1074 652
rect 1355 641 1401 652
rect 1579 793 1625 804
rect 1028 504 1074 606
rect 1579 504 1625 653
rect 1028 458 1484 504
rect 1579 458 1634 504
rect 430 401 534 412
rect 430 355 459 401
rect 505 355 534 401
rect 430 344 534 355
rect 878 401 982 412
rect 878 355 907 401
rect 953 355 982 401
rect 878 344 982 355
rect 1028 264 1074 458
rect 1438 412 1484 458
rect 1214 401 1318 412
rect 1214 355 1243 401
rect 1289 355 1318 401
rect 1214 344 1318 355
rect 1438 401 1542 412
rect 1438 355 1467 401
rect 1513 355 1542 401
rect 1438 344 1542 355
rect 1588 298 1634 458
rect 11 236 1074 264
rect 1579 252 1634 298
rect 57 218 907 236
rect 11 85 57 96
rect 459 142 505 153
rect 459 21 505 96
rect 953 218 1074 236
rect 1355 236 1401 247
rect 907 85 953 96
rect 1355 21 1401 96
rect 1579 237 1625 252
rect 1579 86 1625 97
rect -2 -159 1414 21
<< labels >>
flabel metal1 430 344 534 412 1 FreeSans 192 0 0 0 A
port 1 n
flabel metal1 878 344 982 412 1 FreeSans 192 0 0 0 B
port 2 n
flabel metal1 242 924 316 980 1 FreeSans 192 0 0 0 VDD
port 5 n
flabel nwell -104 706 -30 762 1 FreeSans 192 0 0 0 VNW
port 6 n
flabel pwell -104 76 -30 132 1 FreeSans 192 0 0 0 VPW
port 7 n
flabel metal1 238 -116 312 -60 1 FreeSans 192 0 0 0 VSS
port 8 n
flabel metal1 1243 355 1289 401 1 FreeSans 96 0 0 0 C
port 3 n
flabel metal1 1588 355 1634 401 1 FreeSans 96 0 0 0 Y
port 4 n
flabel metal1 1041 465 1081 495 1 FreeSans 96 0 0 0 idk
<< end >>
