.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.param sw_stat_mismatch=0
.param fnoicor=0
.include maj3.spice
XM0 A B C Y VDD VNW VPW GND maj3
V1 VDD GND 3.3
V2 VNW VDD 0
V3 VPW GND 0
V4 A GND PULSE(0 3.3 0 10p 10p 10n 20n)
V5 B GND PULSE(0 3.3 0 10p 10p 20n 40n)
V6 C GND PULSE(0 3.3 0 10p 10p 40n 80n)
.tran 1p 100n

.control
run
plot v(xm0.idk)+10.5 v(a)-3.5 v(b) v(c)+3.5 v(y)+7
*plot v(a)-3.5 v(b) v(c)+3.5 v(y)+7
.endc
