** sch_path: /foss/designs/real/inyeon-4-chipaton-2025/lvs/gf180mcu_osu_sc_gp9t3v3__maj3.sch
.subckt gf180mcu_osu_sc_gp9t3v3__maj3 VDD VSS A B C Y
*.PININFO VDD:B VSS:B A:I B:I C:I Y:O
M1 net1 C VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M2 X B net1 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M3 net6 A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M5 net2 A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M6 X C net2 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M4 X B net6 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M7 X B net5 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M8 net5 C VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M9 X B net4 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M10 net4 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M11 X C net3 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M12 net3 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M13 Y X VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M14 Y X VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M15 Y X VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M16 Y X VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
.ends
